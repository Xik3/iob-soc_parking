	// SEG
	//input [`SEG_INPUT_W-1:0] seg_input,
	output [3:0] 	seg_anode,   
	output [6:0]    seg_cat,
	output [`SEG_OUTPUT_W-1:0] seg_data_enable,
